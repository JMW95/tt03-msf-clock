module tb (
    input        clk_i,
    input        rst_i,

    input        inc_i,
    output       ovf_o,

    output [1:0] digit_hour_h_o,
    output [3:0] digit_hour_l_o,
    output [2:0] digit_min_h_o,
    output [3:0] digit_min_l_o,
    output [2:0] digit_sec_h_o,
    output [3:0] digit_sec_l_o,

    input        load_i,
    input  [1:0] load_hour_h_i,
    input  [3:0] load_hour_l_i,
    input  [2:0] load_min_h_i,
    input  [3:0] load_min_l_i,
    input  [2:0] load_sec_h_i,
    input  [3:0] load_sec_l_i
);

`ifdef __ICARUS__
    initial begin
        $dumpfile ("tb.vcd");
        $dumpvars (0, tb);
        #1;
    end
`endif

wire hour_l_ovf;
wire min_h_ovf;
wire min_l_ovf;
wire sec_h_ovf;
wire sec_l_ovf;

wire hour_h_at_max;

// 2-bits
digit #(.MAX(2)) hour_h (
    .clk_i        (clk_i),
    .rst_i        (rst_i),
    .digit_o      (digit_hour_h_o),
    .at_max_o     (hour_h_at_max),
    .at_max_i     (1'b0),
    .inc_i        (hour_l_ovf),
    .ovf_o        (ovf_o),
    .load_i       (load_i),
    .load_value_i (load_hour_h_i)
);

// 4-bits
digit #(.MAX(9), .MAX2(3)) hour_l (
    .clk_i        (clk_i),
    .rst_i        (rst_i),
    .digit_o      (digit_hour_l_o),
    .at_max_o     (),
    .at_max_i     (hour_h_at_max),
    .inc_i        (min_h_ovf),
    .ovf_o        (hour_l_ovf),
    .load_i       (load_i),
    .load_value_i (load_hour_l_i)
);

// 3-bits
digit #(.MAX(5)) min_h (
    .clk_i        (clk_i),
    .rst_i        (rst_i),
    .digit_o      (digit_min_h_o),
    .at_max_o     (),
    .at_max_i     (1'b0),
    .inc_i        (min_l_ovf),
    .ovf_o        (min_h_ovf),
    .load_i       (load_i),
    .load_value_i (load_min_h_i)
);

// 4-bits
digit #(.MAX(9)) min_l (
    .clk_i        (clk_i),
    .rst_i        (rst_i),
    .digit_o      (digit_min_l_o),
    .at_max_o     (),
    .at_max_i     (1'b0),
    .inc_i        (sec_h_ovf),
    .ovf_o        (min_l_ovf),
    .load_i       (load_i),
    .load_value_i (load_min_l_i)
);

// 3-bits
digit #(.MAX(5)) sec_h (
    .clk_i        (clk_i),
    .rst_i        (rst_i),
    .digit_o      (digit_sec_h_o),
    .at_max_o     (),
    .at_max_i     (1'b0),
    .inc_i        (sec_l_ovf),
    .ovf_o        (sec_h_ovf),
    .load_i       (load_i),
    .load_value_i (load_sec_h_i)
);

// 4-bits
digit #(.MAX(9)) sec_l (
    .clk_i        (clk_i),
    .rst_i        (rst_i),
    .digit_o      (digit_sec_l_o),
    .at_max_o     (),
    .at_max_i     (1'b0),
    .inc_i        (inc_i),
    .ovf_o        (sec_l_ovf),
    .load_i       (load_i),
    .load_value_i (load_sec_l_i)
);

endmodule
